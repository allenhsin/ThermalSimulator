
module INV_X1M_A12TR
(
    input wire A,
    output wire Y
);

endmodule

module INV_X2M_A12TR (
    Input,
    Output
);

endmodule

module AND_X1M_A12TR ();

    parameter CadenceSucks = 2;
    
endmodule
